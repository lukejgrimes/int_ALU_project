module 4b_and_gate ( input [3:0] a, b, output [3:0] out );
    assign b = a & b;
    
endmodule