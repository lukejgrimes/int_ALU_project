module 4b_div ();

endmodule