module _4b_not_gate( input [3:0] in, output [3:0] out );
    assign out = ~in;
endmodule