module 4b_add ();
    
endmodule