module _2x4_shift (
    input [3:0] a, b,
    
);

endmodule