module 4b_nor_gate(
    input a = 3;
    input b = 0;
    output = y;
);
    assign y = ~(a | b);
endmodule;
