module 4b_mult ();

endmodule