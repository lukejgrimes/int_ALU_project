module 4b_sub ();
    
endmodule